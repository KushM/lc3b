library verilog;
use verilog.vl_types.all;
entity testbenchcontrol is
end testbenchcontrol;
