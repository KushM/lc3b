library verilog;
use verilog.vl_types.all;
entity lc3b is
    port(
        clock           : in     vl_logic;
        reset1          : in     vl_logic
    );
end lc3b;
